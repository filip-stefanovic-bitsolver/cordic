module cordic(
 input clk,
 input rst_n,
 input signed  [15:0] z_tgt,
 output signed [15:0] x_out,
 output signed [15:0] y_out
);
localparam signed[239:0] atan = {16'd1,16'd3,16'd5,16'd10,16'd20,16'd41,16'd81,16'd163,16'd326,16'd652,16'd1302,16'd2594,16'd5110,16'd9672,16'd16384};
reg signed[15:0][15:0] x;
reg signed[15:0][15:0] y;
reg signed[15:0][15:0] z;
reg signed[15:0] z_tmp;
 
always @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    x <= '0;
    y <= '0;
    z <= '0;
  end else begin
    y[0] <= '0;
    z[0] <= z_tgt;
    x[0] <= 16'd19898;
    x[1] <= (!z[0][15]) ? x[0] - (y[0]>>>0) : x[0] + (y[0]>>>0);
    y[1] <= (!z[0][15]) ? y[0] + (x[0]>>>0) : y[0] - (x[0]>>>0);
    z[1] <= (!z[0][15]) ? z[0] - atan[15:0] : z[0] + atan[15:0];
    x[2] <= (!z[1][15]) ? x[1] - (y[1]>>>1) : x[1] + (y[1]>>>1);
    y[2] <= (!z[1][15]) ? y[1] + (x[1]>>>1) : y[1] - (x[1]>>>1);
    z[2] <= (!z[1][15]) ? z[1] - atan[31:16] : z[1] + atan[31:16];
    x[3] <= (!z[2][15]) ? x[2] - (y[2]>>>2) : x[2] + (y[2]>>>2);
    y[3] <= (!z[2][15]) ? y[2] + (x[2]>>>2) : y[2] - (x[2]>>>2);
    z[3] <= (!z[2][15]) ? z[2] - atan[47:32] : z[2] + atan[47:32];
    x[4] <= (!z[3][15]) ? x[3] - (y[3]>>>3) : x[3] + (y[3]>>>3);
    y[4] <= (!z[3][15]) ? y[3] + (x[3]>>>3) : y[3] - (x[3]>>>3);
    z[4] <= (!z[3][15]) ? z[3] - atan[63:48] : z[3] + atan[63:48];
    x[5] <= (!z[4][15]) ? x[4] - (y[4]>>>4) : x[4] + (y[4]>>>4);
    y[5] <= (!z[4][15]) ? y[4] + (x[4]>>>4) : y[4] - (x[4]>>>4);
    z[5] <= (!z[4][15]) ? z[4] - atan[79:64] : z[4] + atan[79:64];
    x[6] <= (!z[5][15]) ? x[5] - (y[5]>>>5) : x[5] + (y[5]>>>5);
    y[6] <= (!z[5][15]) ? y[5] + (x[5]>>>5) : y[5] - (x[5]>>>5);
    z[6] <= (!z[5][15]) ? z[5] - atan[95:80] : z[5] + atan[95:80];
    x[7] <= (!z[6][15]) ? x[6] - (y[6]>>>6) : x[6] + (y[6]>>>6);
    y[7] <= (!z[6][15]) ? y[6] + (x[6]>>>6) : y[6] - (x[6]>>>6);
    z[7] <= (!z[6][15]) ? z[6] - atan[111:96] : z[6] + atan[111:96];
    x[8] <= (!z[7][15]) ? x[7] - (y[7]>>>7) : x[7] + (y[7]>>>7);
    y[8] <= (!z[7][15]) ? y[7] + (x[7]>>>7) : y[7] - (x[7]>>>7);
    z[8] <= (!z[7][15]) ? z[7] - atan[127:112] : z[7] + atan[127:112];
    x[9] <= (!z[8][15]) ? x[8] - (y[8]>>>8) : x[8] + (y[8]>>>8);
    y[9] <= (!z[8][15]) ? y[8] + (x[8]>>>8) : y[8] - (x[8]>>>8);
    z[9] <= (!z[8][15]) ? z[8] - atan[143:128] : z[8] + atan[143:128];
    x[10] <= (!z[9][15]) ? x[9] - (y[9]>>>9) : x[9] + (y[9]>>>9);
    y[10] <= (!z[9][15]) ? y[9] + (x[9]>>>9) : y[9] - (x[9]>>>9);
    z[10] <= (!z[9][15]) ? z[9] - atan[159:144] : z[9] + atan[159:144];
    x[11] <= (!z[10][15]) ? x[10] - (y[10]>>>10) : x[10] + (y[10]>>>10);
    y[11] <= (!z[10][15]) ? y[10] + (x[10]>>>10) : y[10] - (x[10]>>>10);
    z[11] <= (!z[10][15]) ? z[10] - atan[175:160] : z[10] + atan[175:160];
    x[12] <= (!z[11][15]) ? x[11] - (y[11]>>>11) : x[11] + (y[11]>>>11);
    y[12] <= (!z[11][15]) ? y[11] + (x[11]>>>11) : y[11] - (x[11]>>>11);
    z[12] <= (!z[11][15]) ? z[11] - atan[191:176] : z[11] + atan[191:176];
    x[13] <= (!z[12][15]) ? x[12] - (y[12]>>>12) : x[12] + (y[12]>>>12);
    y[13] <= (!z[12][15]) ? y[12] + (x[12]>>>12) : y[12] - (x[12]>>>12);
    z[13] <= (!z[12][15]) ? z[12] - atan[207:192] : z[12] + atan[207:192];
    x[14] <= (!z[13][15]) ? x[13] - (y[13]>>>13) : x[13] + (y[13]>>>13);
    y[14] <= (!z[13][15]) ? y[13] + (x[13]>>>13) : y[13] - (x[13]>>>13);
    z[14] <= (!z[13][15]) ? z[13] - atan[223:208] : z[13] + atan[223:208];
    x[15] <= (!z[14][15]) ? x[14] - (y[14]>>>14) : x[14] + (y[14]>>>14);
    y[15] <= (!z[14][15]) ? y[14] + (x[14]>>>14) : y[14] - (x[14]>>>14);
    z[15] <= (!z[14][15]) ? z[14] - atan[239:224] : z[14] + atan[239:224];
 end
end
assign x_out = (x[15][15] != 1'b1) ? x[15] : 16'd32767;
assign y_out = (y[15][15] != 1'b1) ? y[15] : 16'd32767;
endmodule