module cordic(
 input clk,
 input rst_n,
 input signed  [10:0] z_tgt,
 output signed [10:0] x_out,
 output signed [10:0] y_out
);
localparam signed[109:0] atan = {11'd1,11'd3,11'd5,11'd10,11'd20,11'd41,11'd81,11'd160,11'd302,11'd512};
reg signed[10:0][10:0] x;
reg signed[10:0][10:0] y;
reg signed[10:0][10:0] z;
 
always @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    x <= '0;
    y <= '0;
    z <= '0;
  end else begin
    y[0] <= '0;
    z[0] <= z_tgt;
    x[0] <= 11'd621;
    x[1] <= (!z[0][10]) ? x[0] - (y[0]>>>0) : x[0] + (y[0]>>>0);
    y[1] <= (!z[0][10]) ? y[0] + (x[0]>>>0) : y[0] - (x[0]>>>0);
    z[1] <= (!z[0][10]) ? z[0] - atan[10:0] : z[0] + atan[10:0];
    x[2] <= (!z[1][10]) ? x[1] - (y[1]>>>1) : x[1] + (y[1]>>>1);
    y[2] <= (!z[1][10]) ? y[1] + (x[1]>>>1) : y[1] - (x[1]>>>1);
    z[2] <= (!z[1][10]) ? z[1] - atan[21:11] : z[1] + atan[21:11];
    x[3] <= (!z[2][10]) ? x[2] - (y[2]>>>2) : x[2] + (y[2]>>>2);
    y[3] <= (!z[2][10]) ? y[2] + (x[2]>>>2) : y[2] - (x[2]>>>2);
    z[3] <= (!z[2][10]) ? z[2] - atan[32:22] : z[2] + atan[32:22];
    x[4] <= (!z[3][10]) ? x[3] - (y[3]>>>3) : x[3] + (y[3]>>>3);
    y[4] <= (!z[3][10]) ? y[3] + (x[3]>>>3) : y[3] - (x[3]>>>3);
    z[4] <= (!z[3][10]) ? z[3] - atan[43:33] : z[3] + atan[43:33];
    x[5] <= (!z[4][10]) ? x[4] - (y[4]>>>4) : x[4] + (y[4]>>>4);
    y[5] <= (!z[4][10]) ? y[4] + (x[4]>>>4) : y[4] - (x[4]>>>4);
    z[5] <= (!z[4][10]) ? z[4] - atan[54:44] : z[4] + atan[54:44];
    x[6] <= (!z[5][10]) ? x[5] - (y[5]>>>5) : x[5] + (y[5]>>>5);
    y[6] <= (!z[5][10]) ? y[5] + (x[5]>>>5) : y[5] - (x[5]>>>5);
    z[6] <= (!z[5][10]) ? z[5] - atan[65:55] : z[5] + atan[65:55];
    x[7] <= (!z[6][10]) ? x[6] - (y[6]>>>6) : x[6] + (y[6]>>>6);
    y[7] <= (!z[6][10]) ? y[6] + (x[6]>>>6) : y[6] - (x[6]>>>6);
    z[7] <= (!z[6][10]) ? z[6] - atan[76:66] : z[6] + atan[76:66];
    x[8] <= (!z[7][10]) ? x[7] - (y[7]>>>7) : x[7] + (y[7]>>>7);
    y[8] <= (!z[7][10]) ? y[7] + (x[7]>>>7) : y[7] - (x[7]>>>7);
    z[8] <= (!z[7][10]) ? z[7] - atan[87:77] : z[7] + atan[87:77];
    x[9] <= (!z[8][10]) ? x[8] - (y[8]>>>8) : x[8] + (y[8]>>>8);
    y[9] <= (!z[8][10]) ? y[8] + (x[8]>>>8) : y[8] - (x[8]>>>8);
    z[9] <= (!z[8][10]) ? z[8] - atan[98:88] : z[8] + atan[98:88];
    x[10] <= (!z[9][10]) ? x[9] - (y[9]>>>9) : x[9] + (y[9]>>>9);
    y[10] <= (!z[9][10]) ? y[9] + (x[9]>>>9) : y[9] - (x[9]>>>9);
    z[10] <= (!z[9][10]) ? z[9] - atan[109:99] : z[9] + atan[109:99];
 end
end
assign x_out = x[10];
assign y_out = y[10];
endmodule